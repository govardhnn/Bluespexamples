package clock;

interface Ifc_clock 
(*synthesize*)
module
   
endmodule 
endpackage
