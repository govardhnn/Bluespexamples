function ha(a, b);
   s = a ^ b;
   c = a & b;
   return {c, s};
endfunction
