package full_adder_testbench;

import full_adder :: *;
import half_adder :: *;

(*synthesize*)

module mk_full_adder_testbench(Empty);

// WORK IN PROGRESS


endmodule

endpackage
